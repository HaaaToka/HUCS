module counter(mode, reset, clk, count);
	input mode, reset, clk;
	output[4:0] count;
endmodule
