module four_bit_adder(
    input [3:0] A,
    input [3:0] B,
    input CIN,
    output [4:0] S,
    output COUT
    );

endmodule
